// mymodule.v
module mymodule

// para exportar una funcion tenemos que usar 'pub'
pub fn say_hi() {
	println('Hola desde myfunction...')
}